module priority_encoder_256b(input wire[255:0] in, output reg[7:0] out);
    task encoder_8b (input wire[7:0] dec, output wire[2:0] enc);
    begin
        
    end

    always @* begin
        
    end
endmodule