module core (input clk);

endmodule