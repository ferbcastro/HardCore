module core_TB ();
    reg reset, clk;
    reg[511:0] linha_cache;
    reg[1:0] endereco;

    core DUT(.linha_cache(linha_cache), .endereco(endereco), .clk(clk), .reset(reset));

    initial begin
        // Carrega primeira matriz de assinaturas '[HASH][CLUSTER]'
        $readmemh("./memory_files/primeira_matriz.mem", DUT.primeira_matriz);
        // Carrega segunda matriz de assinaturas '[CLUSTER][HASH]'
        $readmemh("./memory_files/segunda_matriz.mem", DUT.segunda_matriz);
        $dumpfile("core_TB.vcd");
        $dumpvars(2, DUT);
    end

    always #5 clk = ~clk;

    initial begin : BLOCO
        integer i;

        clk = 1'b0;
        reset = 1'b1;
        #1 clk = 1'b1;
        #1 reset = 1'b0;
        clk = 1'b0;
        
        // Colide na hash de XOR mas nao na de ADD
        linha_cache = 512'b00000000001010011110010111001011011011001011100001000000101111010001111000001100100011111111010111010000111011011111100000010101100101011010010001111010001001000101100000110100011101010001101100100110011010010011110111111001010011101010101100000011000000010101101111111100111001010011001101000010011111111010111100101111111001011010011001010110100010100110100101000011100011010000001001100001010101000100110100010100100101011001000101010101010000011000111001001110110001111110100100000001100110001100010000110110;
        endereco = 2'b00;
        #5
        // Malwares codificados nas matrizes
        linha_cache = 512'b01111001001110000110011001000010001001000101110111010111011101001001100001110000000001010000100101010010101000001000011001000111011111110111000101100011011000100010010100101010001000001000010001011100001110011010110001100100110101001011010010100000001010011101001011101111101110011101011111111101100010001000110111000101010111110010010111101101101111110111010011110011000100111010111111000100101011101111100101010000111101110010011011001100101101110100101000101001010110111010100010000011100001011001001010101101;
        endereco = 2'b01;
        #5
        
        for (i = 0; i < 4; i = i + 1) begin
            $display("RESULTADOS[%d] = %d", i, DUT.resultados[i]);
        end

        $stop();
    end
endmodule