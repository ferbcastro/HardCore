module core_TB ();
    reg reset, clk;
    reg[511:0] linha_cache;
    reg[1:0] endereco;

    core DUT(.linha_cache(linha_cache), .endereco(endereco), .clk(clk), .reset(reset));

    initial begin
        // Carrega primeira matriz de assinaturas '[HASH][CLUSTER]'
        $readmemh("./memory_files/primeira_matriz.mem", DUT.primeira_matriz);
        // Carrega segunda matriz de assinaturas '[CLUSTER][HASH]'
        $readmemh("./memory_files/segunda_matriz.mem", DUT.segunda_matriz);
        $dumpfile("core_TB.vcd");
        $dumpvars(2, DUT);
    end

    always #5 clk = ~clk;

    initial begin : BLOCO
        integer i;

        clk = 1'b0;
        reset = 1'b1;
        #1 clk = 1'b1;
        #1 reset = 1'b0;
        clk = 1'b0;
        
        // Colide na hash de XOR mas nao na de ADD
        linha_cache = 512'b00000000001010011110010111001011011011001011100001000000101111010001111000001100100011111111010111010000111011011111100000010101100101011010010001111010001001000101100000110100011101010001101100100110011010010011110111111001010011101010101100000011000000010101101111111100111001010011001101000010011111111010111100101111111001011010011001010110100010100110100101000011100011010000001001100001010101000100110100010100100101011001000101010101010000011000111001001110110001111110100100000001100110001100010000110110;
        endereco = 2'b00;
        #5
        // Malwares codificados nas matrizes
        linha_cache = 512'b00111000011010101110000101110011110100110011101110110101101000101010101001011101000101000010011000101001111011000110011100010000111011011111110000011111011000011000101010011010001110111111111111001111111011110011111000000100100011111000011110001100000001111100000111001110100100010111100100011110100000011111010010100011011100101110001001100011101001101000100010011000011101111011010101000010100111101100110100110010000110011011100010001000001011000100001010000011111110111001110101010101100111100100011111001100;
        endereco = 2'b01;
        #5
        linha_cache = 512'b01001101101110101011011111101000101000100111100011010100010011101001000110100001001000101010111011111010010111000110011001011110001010110110101011100110110100001001100110000101100000000011010000001111011111111011101101010110101000101111000110111000010100000110110011101010011101001010110100100100100011100110100100010010110110100001110101001110011101010000001010101111111110111110001101010110010001010100000101011100001000101110110000001111110101101101110001101100000101010011111110111001001000011110110100101000;
        endereco = 2'b10;
        #5
        
        for (i = 0; i < 4; i = i + 1) begin
            $display("RESULTADOS[%d] = %d", i, DUT.resultados[i]);
        end

        $stop();
    end
endmodule