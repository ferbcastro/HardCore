module core_TB ();

    initial begin
        
    end

    always

    initial begin
        $stop()
    end

endmodule