module xor_hash_TB ();
    reg[511:0] entrada;
    wire[7:0] saida;

    xor_hash DUT(.in(entrada), .out(saida));

    initial begin
        // $monitor("saida = %d", saida);
    end

    initial begin
        // entrada = {511'b0, 1'b1};
        // #5 entrada = {503'b0, 1'b1, 8'b00000001};
           entrada = 512'b11010000001010010000111110001100101111010001100111101100010010100110011101100111010011101111000110111101101100000101000001111100111100110000111101100001000101111000011110001101000111111010110100111110101000111100100010110001100101010000001001110100001000110111111010011111111100100011100110011111110100011011101010101100001011011101001100111110101001010000010001101110001001100110110101111001011110001010101100101100110010100011001110111111011001000101001001010101000111111011011100010101100101110011000110011010;
        #5 $display("saida = %d", saida); entrada = 512'b00111000011010101110000101110011110100110011101110110101101000101010101001011101000101000010011000101001111011000110011100010000111011011111110000011111011000011000101010011010001110111111111111001111111011110011111000000100100011111000011110001100000001111100000111001110100100010111100100011110100000011111010010100011011100101110001001100011101001101000100010011000011101111011010101000010100111101100110100110010000110011011100010001000001011000100001010000011111110111001110101010101100111100100011111001100;
        #5 $display("saida = %d", saida); entrada = 512'b01001101101110101011011111101000101000100111100011010100010011101001000110100001001000101010111011111010010111000110011001011110001010110110101011100110110100001001100110000101100000000011010000001111011111111011101101010110101000101111000110111000010100000110110011101010011101001010110100100100100011100110100100010010110110100001110101001110011101010000001010101111111110111110001101010110010001010100000101011100001000101110110000001111110101101101110001101100000101010011111110111001001000011110110100101000;
        #5 $display("saida = %d", saida); entrada = 512'b10011001000110110101110111110001001011101011110100110100000010000010000110110001011100010110100110011110010010101000011101100010111101110100100100010000110011101110001100100110110100011100100111110010010000000011001111000111000010101100000010100100100001100000110101001000101100000000111110110011100111000010011110110100010111111110001101000101011001010010110111010000001010011010101001111000001010101001111001000000110010100001110100011001011100111011101000011101000111100110001010110011111100011010100110110011; 
        #5 $display("saida = %d", saida); entrada = 512'b01010100101000111011011101010000101111101100011111110101000010000100000000100100000110011101110111100111111100001101110100000001001101100100001100011000001110011101001001010111100000001111001011110011000111101111110010100100111100011000000011010100100010011100000000111110100001001101111010100001001110100111011001110100000001110110010000100010111111100000111101110111101011001110101100011000101001101011101110100000010111100010100111111011000110011110000011011001010110000010001001000011101011001110001001001100; 
        #5 $display("saida = %d", saida); entrada = 512'b10001011001010000000101000111010111010111101101000001001001100011101010001110000000111000000111111111011110001000010011010111010010101010101101110101111111000111011100011001100111010011011001111011110110000000110010100000111010001100011001101001100001111101011001100101110010001111111111000000110111100000000010000111011100101111100011111111001101010000000100000111000100010001111101010111100011010000111011001110011110000100100110111001100101010010011101101111111100111100000000101000100001000110111010001110000; 
        #5 $display("saida = %d", saida); entrada = 512'b10000001001100001100001000011000001011000000110011010101100110011110110010111000001110011110000000011010110001000010110100001001001010000100100110000011101111001101111000110011111100010101001100010111101111001010100100010101010111111100100000000010001100101111111000100001001100101100000100011100101010101101111001010110110110000011001101001011011001001011100111100010000111110011100110000100110011100011111010000010011001111011001100111001100001011001101110101111111000010010011111000100111100100100000011111000; 
        #5 $display("saida = %d", saida); entrada = 512'b01111001001110000110011001000010001001000101110111010111011101001001100001110000000001010000100101010010101000001000011001000111011111110111000101100011011000100010010100101010001000001000010001011100001110011010110001100100110101001011010010100000001010011101001011101111101110011101011111111101100010001000110111000101010111110010010111101101101111110111010011110011000100111010111111000100101011101111100101010000111101110010011011001100101101110100101000101001010110111010100010000011100001011001001010101101;
        #5 $display("saida = %d", saida); entrada = 512'b00000000001010011110010111001011011011001011100001000000101111010001111000001100100011111111010111010000111011011111100000010101100101011010010001111010001001000101100000110100011101010001101100100110011010010011110111111001010011101010101100000011000000010101101111111100111001010011001101000010011111111010111100101111111001011010011001010110100010100110100101000011100011010000001001100001010101000100110100010100100101011001000101010101010000011000111001001110110001111110100100000001100110001100010000110110;
        #5 $display("saida = %d", saida); $finish();
    end
endmodule